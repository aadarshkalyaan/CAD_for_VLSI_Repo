package MAC_Wrapper;
import FIFO::*;
import CAD_V1::*;
import SpecialFIFOs::*;

interface MAC_Wrapper_IFC;
    // Input methods
    method Action enqS(Bit#(1) s);
    method Action enqB(Bit#(16) b);
    method Action enqC(Bit#(32) c);
    method Action enqA(Bit#(16) a);
    
    // Pass-through output methods
    method ActionValue#(Bit#(16)) get_a_out();  
    method ActionValue#(Bit#(16)) get_b_out();  
    method ActionValue#(Bit#(1)) get_s_out();   
    
    // MAC computation output
    method ActionValue#(Bit#(32)) get_MAC_result();
endinterface

(* synthesize *)
module mkMAC_Wrapper(MAC_Wrapper_IFC);
    // Input FIFOs
    FIFO#(Bit#(1)) s_fifo <- mkPipelineFIFO;
    FIFO#(Bit#(16)) b_fifo <- mkPipelineFIFO;
    FIFO#(Bit#(32)) c_fifo <- mkPipelineFIFO;
    FIFO#(Bit#(16)) a_fifo <- mkPipelineFIFO;
    
    // Output FIFOs for pass-through
    FIFO#(Bit#(16)) a_out_fifo <- mkPipelineFIFO;
    FIFO#(Bit#(16)) b_out_fifo <- mkPipelineFIFO;
    FIFO#(Bit#(1)) s_out_fifo <- mkPipelineFIFO;
    
    // Output FIFO for MAC result
    FIFO#(Bit#(32)) mac_result_fifo <- mkPipelineFIFO;
    
    // Instantiate the MAC module
    TOP_IFC mac <- mkMAC();
    
    // Rule to handle pass-through and MAC computation
    rule process_inputs;
        let s = s_fifo.first;
        let b = b_fifo.first;
        let c = c_fifo.first;
        let a = a_fifo.first;
        
        // Compute MAC result
        let mac_result = mac.get_MAC(a, b, c, s);
        
        // Enqueue to output FIFOs
        a_out_fifo.enq(a);
        b_out_fifo.enq(b);
        s_out_fifo.enq(s);
        mac_result_fifo.enq(mac_result);
        
        // Dequeue from input FIFOs
        s_fifo.deq;
        b_fifo.deq;
        c_fifo.deq;
        a_fifo.deq;
    endrule
    
    // Input methods
    method Action enqS(Bit#(1) s);
        s_fifo.enq(s);
    endmethod
    
    method Action enqB(Bit#(16) b);
        b_fifo.enq(b);
    endmethod
    
    method Action enqC(Bit#(32) c);
        c_fifo.enq(c);
    endmethod
    
    method Action enqA(Bit#(16) a);
        a_fifo.enq(a);
    endmethod
    
    // Pass-through output methods
    method ActionValue#(Bit#(16)) get_a_out();
        a_out_fifo.deq;
        return a_out_fifo.first;
    endmethod
    
    method ActionValue#(Bit#(16)) get_b_out();
        b_out_fifo.deq;
        return b_out_fifo.first;
    endmethod
    
    method ActionValue#(Bit#(1)) get_s_out();
        s_out_fifo.deq;
        return s_out_fifo.first;
    endmethod
    
    // MAC result output method
    method ActionValue#(Bit#(32)) get_MAC_result();
        mac_result_fifo.deq;
        return mac_result_fifo.first;
    endmethod
endmodule

endpackage