package rca;
    interface Action start(Bit#(32) a,)
endpackage;